module mux4(ALUSel_reg);
output reg [2:0] ALUSel_reg;
endmodule